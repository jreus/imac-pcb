* NXP Semiconductors
.subckt PemiQFN_HT INPUT1 PADGND OUTPUT1
C1  1   500 .053p
C2  2   500 .053p
C3  3   500 .053p
C4  4   500 .053p
C5  5   500 .053p
C6  6   500 .053p
C7  7   500 .053p
C8  8   500 .053p
C9  9   500 .053p
C10 10  500 .053p
C11 11  500 .053p
C12 12  500 .053p
C13 13  500 .053p
C14 14  500 .053p
C15 15  500 .053p
C16 16  500 .053p
C17 17  500 .053p
C18 18  500 .053p
C19 19  500 .053p
R1  1  2  2.250
R2  2  3  2.250
R3  3  4  2.250
R4  4  5  2.250
R5  5  6  2.250
R6  6  7  2.250
R7  7  8  2.250
R8  8  9  2.250
R9  9  10 2.250
R10 10 11 2.250
R11 11 12 2.250
R12 12 13 2.250
R13 13 14 2.250
R14 14 15 2.250
R15 15 16 2.250
R16 16 17 2.250
R17 17 18 2.250
R18 18 19 2.250
R19 19 201 2.250
R20 1  101 2.250
D1  500 101 IDS_diode
D2  500 201 IDS_diode
L1  INPUT1  100  400p
L2  OUTPUT1 200  400p
L3  500   501    25p
R200 201  200    0.020
R100 100  101    0.020
R300 501  PADGND 0.2
.model IDS_diode D (VJ = 600m BV = 8 CJO = 19.500p M = 360m)
.ends PemiQFN_HT
