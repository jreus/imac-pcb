* NXP Semiconductors
.subckt PemiQFN_WK INPUT1 PADGND OUTPUT1
C1  1   500 .053p
C2  2   500 .053p
C3  3   500 .053p
C4  4   500 .053p
C5  5   500 .053p
C6  6   500 .053p
C7  7   500 .053p
C8  8   500 .053p
C9  9   500 .053p
C10 10  500 .053p
C11 11  500 .053p
C12 12  500 .053p
C13 13  500 .053p
C14 14  500 .053p
C15 15  500 .053p
C16 16  500 .053p
C17 17  500 .053p
C18 18  500 .053p
C19 19  500 .053p
R1  1  2  10.000
R2  2  3  10.000
R3  3  4  10.000
R4  4  5  10.000
R5  5  6  10.000
R6  6  7  10.000
R7  7  8  10.000
R8  8  9  10.000
R9  9  10 10.000
R10 10 11 10.000
R11 11 12 10.000
R12 12 13 10.000
R13 13 14 10.000
R14 14 15 10.000
R15 15 16 10.000
R16 16 17 10.000
R17 17 18 10.000
R18 18 19 10.000
R19 19 201 10.000
R20 1  101 10.000
D1  500 101 IDS_diode
D2  500 201 IDS_diode
L1  INPUT1  100  400p
L2  OUTPUT1 200  400p
L3  500   501    25p
R200 201  200    0.020
R100 100  101    0.020
R300 501  PADGND 0.2
.model IDS_diode D (VJ = 600m BV = 8 CJO = 11.000p M = 360m)
.ends PemiQFN_WK
